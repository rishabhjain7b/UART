// Transmitter module for UART


