// 8 bit counter for Baud Rate Generator of UART

module counter_8bit #(parameter limit = 2)
(input clkdiv,
 output reg out);

reg [7:0]k=8'd0;

always @ (posedge clkdiv)
begin
	if (k == (limit-1))
	begin
		k <= 0;
		out <= 0;
	end
	else
	begin
		k <= k+1;
		out <= 1;
	end
end
endmodule

