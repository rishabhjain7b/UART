// Transmitter module for UART

module uart_tx #(parameter data_bits=8, parameter transmitted_bit_counter_bits=4, parameter br=3'b000)
(input [data_bits-1:0]DBUS,
 input sysclk,rst_n,txd_startH,
 output txd,txd_doneH);

 wire bclk;
 wire shftTSR,loadTSR,start;
 wire clr,inc;
 wire [transmitted_bit_counter_bits-1:0]bct;
 wire txd_done,bclk_dlayed;
 wire bclk_rising;

 BRG #(.sel(br)) baud_rate_generator (.fclk(sysclk),.bclkx8(),.bclk(bclk));

 dff DFF1 (.clk(sysclk),.rst_n(rst_n),.in(bclk),.q(bclk_dlayed));
 
 and and_gate (bclk_rising,bclk,~(bclk_dlayed));
 
 sm_tx #(.data_bits(data_bits)) state_machine (.bclk(bclk_rising),.rst_n(rst_n),.txd_startH(txd_startH),.bct(bct),
 						.txd_done(txd_done),.start(start),.shftTSR(shftTSR),.loadTSR(loadTSR),
						.clr(clr),.inc(inc));

 counter_nbit #(.n(transmitted_bit_counter_bits)) transmitted_bit_counter (.clk(sysclk),.clear(clr),.inc(inc),.out(bct));

 PISO #(.piso_width(data_bits)) data_shift_register (.clk(sysclk),.shift(shftTSR),.start(start),.load(loadTSR),.in(DBUS),.out(txd));

 dff DFF2 (.clk(sysclk),.rst_n(rst_n),.in(txd_done),.q(txd_doneH));

endmodule
